module main

import vmir

fn main() {
	
}