module test

import vmir



pub fn test_output() {
}

pub fn test_scan_string() {
}

pub fn test_write() {
}

pub fn test_read() {
}

pub fn test_write_with_func() {
}

pub fn test_read_with_func() {
}
