module test

import vmir

pub fn test_init_context() {
	
	assert true
}