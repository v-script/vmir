module vmir

// context
fn init_context() {
}

fn finist_context() {
}

fn output() {
}

fn scan_string() {
}

fn write() {
}

fn write_with_func() {
}

fn read() {
}

fn read_with_func() {
}

// module
fn new_module() {
}

fn finish_module() {
}

fn get_module_list() {
}

fn new_import() {
}

fn new_export() {
}

fn new_forword() {
}

fn new_proto_arr() {
}

fn new_proto() {
}

fn new_vararg_proto_arr() {
}

fn new_vararg_proto() {
}

// func
fn new_func_arr() {
}

fn new_func() {
}

fn new_vararg_func_arr() {
}

fn new_vararg_func() {
}

fn new_func_reg() {
}

fn finish_func() {
}

fn new_data() {
}

fn new_string_data() {
}

fn new_ref_data() {
}

fn new_expr_data() {
}

fn new_bss() {
}

fn output_item() {
}

fn output_module() {
}

// operands

fn new_int_op() {
}

fn new_uint_op() {
}

fn new_float_op() {
}

fn new_double_op() {
}

fn new_ldouble_op() {
}

fn new_str_op() {
}

fn new_label() {
}

fn new_ref_op() {
}

fn new_reg_op() {
}

fn new_mem_op() {
}

fn output_op() {
}

// insn
fn new_insn() {
}

fn new_insn_arr() {
}

fn new_call_insn() {
}

fn new_ret_insn() {
}

fn prepend_insn() {
}

fn append_insn() {
}

fn insert_insn_after() {
}

fn insert_insn_before() {
}

fn remove_insn() {
}

fn output_insn() {
}

// other api
fn get_error_func() {
}

fn set_error_func() {
}

fn load_module() {
}

fn load_external() {
}

fn link() {
}

// run with interpreter
fn interp() {
}

fn set_interp_interface() {
}

// generator
fn gen_init() {
}

fn gen_finish() {
}

fn gen() {
}

fn set_degug_file() {
}

fn gen_set_debug_level() {
}

fn gen_set_optimize_level() {
}
