module vmir

